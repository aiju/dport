`timescale 1 ns / 1 ps
`default_nettype none

`define ATTRMAX 208
`define symBS 8'hbc
`define symBE 8'hfb
`define symSS 8'h5c
`define symSE 8'hfd
`define symFS 8'hfe
`define symFE 8'hf7
`define symSR 8'h1c
